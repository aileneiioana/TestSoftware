
module hw_nios (
	clk_clk,
	reset_reset_n,
	pio_0_external_connection_export);	

	input		clk_clk;
	input		reset_reset_n;
	output		pio_0_external_connection_export;
endmodule
